//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: FPGA Verilog full testbench for top-level netlist of design: and2_latch
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Wed Aug 16 14:34:16 2023
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

//----- Default net type -----
`default_nettype none

module and2_latch_autocheck_top_tb;
// ----- Local wires for global ports of FPGA fabric -----
wire [0:0] set;
wire [0:0] reset;
wire [0:0] clk;

// ----- Local wires for I/Os of FPGA fabric -----
wire [0:31] gfpga_pad_GPIO_PAD;



reg [0:0] __config_done__;
wire [0:0] __prog_clock__;
reg [0:0] __prog_clock___reg__;
wire [0:0] __op_clock__;
reg [0:0] __op_clock___reg__;
reg [0:0] __prog_reset__;
reg [0:0] __prog_set_;
reg [0:0] __greset__;
reg [0:0] __gset__;
// ---- Address port for Bit-Line decoder -----
reg [0:4] bl_address;
// ---- Address port for Word-Line decoder -----
reg [0:4] wl_address;
// ---- Data input port for memory decoders -----
reg [0:0] data_in;
// ---- Readback port for memory decoders -----
// ---- Wire enable port of memory decoders  -----
wire [0:0] enable;
reg [0:0] enable_reg__;
	assign enable[0]= ~enable_reg__[0] & ~__config_done__[0];
// ----- Shared inputs -------
	reg [0:0] a_shared_input;
	reg [0:0] b_shared_input;

// ----- FPGA fabric outputs -------
	wire [0:0] c_fpga;
	wire [0:0] d_fpga;

// ----- Benchmark outputs -------
	wire [0:0] c_benchmark;
	wire [0:0] d_benchmark;

// ----- Output vectors checking flags -------
	reg [0:0] c_flag;
	reg [0:0] d_flag;

// ----- Error counter: Deposit an error for config_done signal is not raised at the beginning -----
	integer nb_error= 1;
// ----- Number of clock cycles in configuration phase: 615 -----
// ----- Begin configuration done signal generation -----
initial
	begin
		__config_done__[0] = 1'b0;
	end

// ----- End configuration done signal generation -----

// ----- Begin raw programming clock signal generation -----
initial
	begin
		__prog_clock___reg__[0] = 1'b0;
	end
always
	begin
		#5	__prog_clock___reg__[0] = ~__prog_clock___reg__[0];
	end

// ----- End raw programming clock signal generation -----

// ----- Actual programming clock is triggered only when __config_done__ and __prog_reset__ are disabled -----
	assign __prog_clock__[0] = __prog_clock___reg__[0] & (~__config_done__[0]) & (~__prog_reset__[0]);

// ----- Begin raw operating clock signal generation -----
initial
	begin
		__op_clock___reg__[0] = 1'b0;
	end
always wait(~__greset__)
	begin
		#0.4702859819	__op_clock___reg__[0] = ~__op_clock___reg__[0];
	end

// ----- End raw operating clock signal generation -----
// ----- Actual operating clock is triggered only when __config_done__ is enabled -----
	assign __op_clock__[0] = __op_clock___reg__[0] & __config_done__[0];

// ----- Begin programming reset signal generation -----
initial
	begin
		__prog_reset__[0] = 1'b1;
	#10	__prog_reset__[0] = 1'b0;
	end

// ----- End programming reset signal generation -----

// ----- Begin programming set signal generation -----
initial
	begin
		__prog_set_[0] = 1'b1;
	#10	__prog_set_[0] = 1'b0;
	end

// ----- End programming set signal generation -----

// ----- Begin operating reset signal generation -----
// ----- Reset signal is enabled until the first clock cycle in operation phase -----
initial
	begin
		__greset__[0] = 1'b1;
	wait(__config_done__)
	#0.9405719638	__greset__[0] = 1'b1;
	#1.881143928	__greset__[0] = 1'b0;
	end

// ----- End operating reset signal generation -----
// ----- Begin operating set signal generation: always disabled -----
initial
	begin
		__gset__[0] = 1'b0;
	end

// ----- End operating set signal generation: always disabled -----

// ---- Generate enable signal waveform  -----
initial
	begin
		enable_reg__[0] = 1'b0;
		#2.5;
		forever enable_reg__[0] = #5 ~enable_reg__[0];
	end

// ----- Begin connecting global ports of FPGA fabric to stimuli -----
	assign clk[0] = __op_clock__[0];
	assign reset[0] = __greset__[0];
	assign set[0] = __gset__[0];
// ----- End connecting global ports of FPGA fabric to stimuli -----
// ----- FPGA top-level module to be capsulated -----
	fpga_top FPGA_DUT (
		.set(set[0]),
		.reset(reset[0]),
		.clk(clk[0]),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[0:31]),
		.enable(enable[0]),
		.bl_address(bl_address[0:4]),
		.wl_address(wl_address[0:4]),
		.data_in(data_in[0]));

// ----- Link BLIF Benchmark I/Os to FPGA I/Os -----
// ----- Blif Benchmark input a is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD[15] -----
	assign gfpga_pad_GPIO_PAD[15] = a_shared_input[0];

// ----- Blif Benchmark input b is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD[30] -----
	assign gfpga_pad_GPIO_PAD[30] = b_shared_input[0];

// ----- Blif Benchmark input clk is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD[11] -----
	assign gfpga_pad_GPIO_PAD[11] = clk[0];

// ----- Blif Benchmark output c is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD[12] -----
	assign c_fpga[0] = gfpga_pad_GPIO_PAD[12];

// ----- Blif Benchmark output d is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD[26] -----
	assign d_fpga[0] = gfpga_pad_GPIO_PAD[26];

// ----- Wire unused FPGA I/Os to constants -----
	assign gfpga_pad_GPIO_PAD[0] = 1'b0;
	assign gfpga_pad_GPIO_PAD[1] = 1'b0;
	assign gfpga_pad_GPIO_PAD[2] = 1'b0;
	assign gfpga_pad_GPIO_PAD[3] = 1'b0;
	assign gfpga_pad_GPIO_PAD[4] = 1'b0;
	assign gfpga_pad_GPIO_PAD[5] = 1'b0;
	assign gfpga_pad_GPIO_PAD[6] = 1'b0;
	assign gfpga_pad_GPIO_PAD[7] = 1'b0;
	assign gfpga_pad_GPIO_PAD[8] = 1'b0;
	assign gfpga_pad_GPIO_PAD[9] = 1'b0;
	assign gfpga_pad_GPIO_PAD[10] = 1'b0;
	assign gfpga_pad_GPIO_PAD[13] = 1'b0;
	assign gfpga_pad_GPIO_PAD[14] = 1'b0;
	assign gfpga_pad_GPIO_PAD[16] = 1'b0;
	assign gfpga_pad_GPIO_PAD[17] = 1'b0;
	assign gfpga_pad_GPIO_PAD[18] = 1'b0;
	assign gfpga_pad_GPIO_PAD[19] = 1'b0;
	assign gfpga_pad_GPIO_PAD[20] = 1'b0;
	assign gfpga_pad_GPIO_PAD[21] = 1'b0;
	assign gfpga_pad_GPIO_PAD[22] = 1'b0;
	assign gfpga_pad_GPIO_PAD[23] = 1'b0;
	assign gfpga_pad_GPIO_PAD[24] = 1'b0;
	assign gfpga_pad_GPIO_PAD[25] = 1'b0;
	assign gfpga_pad_GPIO_PAD[27] = 1'b0;
	assign gfpga_pad_GPIO_PAD[28] = 1'b0;
	assign gfpga_pad_GPIO_PAD[29] = 1'b0;
	assign gfpga_pad_GPIO_PAD[31] = 1'b0;

// ----- Reference Benchmark Instanication -------
	and2_latch REF_DUT(
		.a(a_shared_input),
		.b(b_shared_input),
		.clk(clk),
		.c(c_benchmark),
		.d(d_benchmark)
	);
// ----- End reference Benchmark Instanication -------

`define BITSTREAM_LENGTH 614
`define BITSTREAM_WIDTH 11
// ----- Virtual memory to store the bitstream from external file -----
reg [0:`BITSTREAM_WIDTH - 1] bit_mem[0:`BITSTREAM_LENGTH - 1];
reg [$clog2(`BITSTREAM_LENGTH):0] bit_index;
// ----- Preload bitstream file to a virtual memory -----
initial begin
	$readmemb("fabric_bitstream.bit", bit_mem);
// ----- Bit-Line Address port default input -----
	bl_address[0:4] = {5{1'b0}};
// ----- Word-Line Address port default input -----
	wl_address[0:4] = {5{1'b0}};
// ----- Data-input port default input -----
	data_in[0] = 1'b0;
	bit_index <= 0;
end
// ----- Begin bitstream loading during configuration phase -----
always @(negedge __prog_clock___reg__[0]) begin
	if (bit_index >= `BITSTREAM_LENGTH) begin
		__config_done__[0] <= 1'b1;
	end else begin
		{bl_address[0:4], wl_address[0:4], data_in[0]} <= bit_mem[bit_index];
		bit_index <= bit_index + 1;
	end
end
// ----- End bitstream loading during configuration phase -----

// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_3_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_2.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_2.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_2.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_2.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_4.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_4.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_4.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_4.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_6.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_6.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_6.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_6.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_8.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_8.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_8.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_8.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_10.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_10.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_10.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_10.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_12.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_12.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_12.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_12.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_14.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_14.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_14.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_14.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_16.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_16.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_16.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_16.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_2.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_2.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_2.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_2.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_4.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_4.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_4.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_4.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_6.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_6.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_6.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_6.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_8.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_8.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_8.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_8.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_10.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_10.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_10.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_10.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_12.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_12.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_12.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_12.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_14.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_14.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_14.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_14.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_16.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_16.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_16.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_16.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_2.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_2.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_2.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_2.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_4.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_4.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_4.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_4.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_6.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_6.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_6.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_6.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_8.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_8.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_8.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_8.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_10.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_10.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_10.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_10.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_12.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_12.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_12.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_12.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_14.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_14.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_14.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_14.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_16.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_16.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_16.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_16.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_2.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_2.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_2.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_2.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_4.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_4.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_4.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_4.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_6.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_6.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_6.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_6.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_8.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_8.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_8.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_8.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_10.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_10.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_10.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_10.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_12.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_12.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_12.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_12.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_14.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_14.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_14.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_14.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_16.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_16.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_16.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_16.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_3.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_3.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_3.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_3.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_5.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_5.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_5.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_5.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_7.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_7.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_7.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_7.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_9.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_9.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_9.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_9.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_11.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_11.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_11.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_11.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_13.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_13.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_13.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_13.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_15.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_15.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_15.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_15.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_17.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_17.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_17.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_17.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_3.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_3.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_3.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_3.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_5.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_5.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_5.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_5.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_7.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_7.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_7.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_7.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_9.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_9.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_9.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_9.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_11.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_11.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_11.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_11.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_13.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_13.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_13.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_13.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_15.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_15.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_15.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_15.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_17.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_17.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_17.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_17.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_3.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_3.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_3.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_3.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_4.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_4.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_4.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_4.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_5.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_5.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_5.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_5.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_6.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_6.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_6.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_6.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_6.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_7.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_7.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_7.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_2.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_3.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_3.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_3.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_3.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_3.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_4.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_4.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_4.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_4.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_4.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_5.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_5.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_5.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_5.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_6.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_6.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_6.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_6.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_6.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_6.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_7.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_7.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_7.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_7.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_7.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_1.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_1.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_2.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_2.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_2.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_2.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_2.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_2.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_2.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_2.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_2.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_3.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_3.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_3.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_3.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_3.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_3.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_3.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_3.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_4.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_4.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_4.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_4.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_4.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_4.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_4.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_4.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_4.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_5.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_5.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_5.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_5.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_5.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_5.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_5.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_5.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_5.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_6.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_6.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_6.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_6.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_6.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_6.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_6.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_6.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_6.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_7.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_7.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_7.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_7.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_7.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_7.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_7.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_7.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_7.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ----- Begin reset signal generation -----
// ----- Input Initialization -------
	initial begin
		a_shared_input <= 1'b0;
		b_shared_input <= 1'b0;

		c_flag[0] <= 1'b0;
		d_flag[0] <= 1'b0;
	end

// ----- Input Stimulus -------
	always@(negedge __op_clock__[0]) begin
		a_shared_input <= $random;
		b_shared_input <= $random;
	end

// ----- Begin checking output vectors -------
// ----- Skip the first falling edge of clock, it is for initialization -------
	reg [0:0] sim_start;

	always@(negedge clk[0]) begin
		if (1'b1 == sim_start[0]) begin
			sim_start[0] <= ~sim_start[0];
		end else 
if (1'b1 == __config_done__) begin
			if(!(c_fpga === c_benchmark) && !(c_benchmark === 1'bx)) begin
				c_flag <= 1'b1;
			end else begin
				c_flag<= 1'b0;
			end
			if(!(d_fpga === d_benchmark) && !(d_benchmark === 1'bx)) begin
				d_flag <= 1'b1;
			end else begin
				d_flag<= 1'b0;
			end
		end
	end

	always@(posedge c_flag) begin
		if(c_flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on c_fpga at time = %t", $realtime);
		end
	end

	always@(posedge d_flag) begin
		if(d_flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on d_fpga at time = %t", $realtime);
		end
	end


// ----- Configuration done must be raised in the end -------
	always@(posedge __config_done__[0]) begin
		nb_error = nb_error - 1;
	end

// ----- Begin output waveform to VCD file-------
	initial begin
		$dumpfile("and2_latch_formal.vcd");
		$dumpvars(1, and2_latch_autocheck_top_tb);
	end
// ----- END output waveform to VCD file -------

initial begin
	sim_start[0] <= 1'b1;
	$timeformat(-9, 2, "ns", 20);
	$display("Simulation start");
// ----- Can be changed by the user for his/her need -------
	#6174
	if(nb_error == 0) begin
		$display("Simulation Succeed");
	end else begin
		$display("Simulation Failed with %d error(s)", nb_error);
	end
	$finish;
end

endmodule
// ----- END Verilog module for and2_latch_autocheck_top_tb -----

//----- Default net type -----
`default_nettype none


//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for physical tile: clb]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Wed Aug 16 14:34:46 2023
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

// ----- BEGIN Grid Verilog module: grid_clb -----
//----- Default net type -----
`default_nettype none

// ----- Verilog module for grid_clb -----
module grid_clb(set,
                reset,
                clk,
                top_width_0_height_0_subtile_0__pin_I_0_,
                top_width_0_height_0_subtile_0__pin_I_4_,
                top_width_0_height_0_subtile_0__pin_I_8_,
                right_width_0_height_0_subtile_0__pin_I_1_,
                right_width_0_height_0_subtile_0__pin_I_5_,
                right_width_0_height_0_subtile_0__pin_I_9_,
                bottom_width_0_height_0_subtile_0__pin_I_2_,
                bottom_width_0_height_0_subtile_0__pin_I_6_,
                bottom_width_0_height_0_subtile_0__pin_clk_0_,
                left_width_0_height_0_subtile_0__pin_I_3_,
                left_width_0_height_0_subtile_0__pin_I_7_,
                bl,
                wl,
                top_width_0_height_0_subtile_0__pin_O_2_,
                right_width_0_height_0_subtile_0__pin_O_3_,
                bottom_width_0_height_0_subtile_0__pin_O_0_,
                left_width_0_height_0_subtile_0__pin_O_1_);
//----- GLOBAL PORTS -----
input [0:0] set;
//----- GLOBAL PORTS -----
input [0:0] reset;
//----- GLOBAL PORTS -----
input [0:0] clk;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I_4_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_I_8_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_I_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_I_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_I_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_I_3_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_I_7_;
//----- INPUT PORTS -----
input [0:14] bl;
//----- INPUT PORTS -----
input [0:13] wl;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_O_2_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_O_3_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_O_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_O_1_;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	logical_tile_clb_mode_clb_ logical_tile_clb_mode_clb__0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.clb_I({top_width_0_height_0_subtile_0__pin_I_0_, right_width_0_height_0_subtile_0__pin_I_1_, bottom_width_0_height_0_subtile_0__pin_I_2_, left_width_0_height_0_subtile_0__pin_I_3_, top_width_0_height_0_subtile_0__pin_I_4_, right_width_0_height_0_subtile_0__pin_I_5_, bottom_width_0_height_0_subtile_0__pin_I_6_, left_width_0_height_0_subtile_0__pin_I_7_, top_width_0_height_0_subtile_0__pin_I_8_, right_width_0_height_0_subtile_0__pin_I_9_}),
		.clb_clk(bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.bl({bl[0:14], bl[0:14], bl[0:14], bl[0:14], bl[0:14], bl[0:14], bl[0:14], bl[0:14], bl[0:14], bl[0:14], bl[0:14], bl[0:14], bl[0:14], bl[0:8]}),
		.wl({wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0], wl[0:1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1], wl[1:2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2], wl[2:3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3], wl[3:4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4], wl[4:5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5], wl[5:6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6], wl[6:7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7], wl[7:8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8], wl[8:9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9], wl[9:10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10], wl[10:11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11], wl[11:12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12], wl[12:13], wl[13], wl[13], wl[13], wl[13], wl[13], wl[13], wl[13], wl[13]}),
		.clb_O({bottom_width_0_height_0_subtile_0__pin_O_0_, left_width_0_height_0_subtile_0__pin_O_1_, top_width_0_height_0_subtile_0__pin_O_2_, right_width_0_height_0_subtile_0__pin_O_3_}));

endmodule
// ----- END Verilog module for grid_clb -----

//----- Default net type -----
`default_nettype none



// ----- END Grid Verilog module: grid_clb -----


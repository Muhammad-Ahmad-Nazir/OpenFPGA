//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: FPGA Verilog full testbench for top-level netlist of design: or2
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Wed Aug 16 11:44:21 2023
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

//----- Default net type -----
`default_nettype none

module or2_autocheck_top_tb;
// ----- Local wires for global ports of FPGA fabric -----
wire [0:0] prog_clk;
wire [0:0] set;
wire [0:0] reset;
wire [0:0] clk;

// ----- Local wires for I/Os of FPGA fabric -----
wire [0:31] gfpga_pad_GPIO_PAD;



reg [0:0] __config_done__;
wire [0:0] __prog_clock__;
reg [0:0] __prog_clock___reg__;
wire [0:0] __op_clock__;
reg [0:0] __op_clock___reg__;
reg [0:0] __prog_reset__;
reg [0:0] __prog_set_;
reg [0:0] __greset__;
reg [0:0] __gset__;
// ---- Configuration-chain head -----
reg [0:0] ccff_head;
// ---- Configuration-chain tail -----
wire [0:0] ccff_tail;
// ----- Shared inputs -------
	reg [0:0] a_shared_input;
	reg [0:0] b_shared_input;

// ----- FPGA fabric outputs -------
	wire [0:0] c_fpga;

// ----- Benchmark outputs -------
	wire [0:0] c_benchmark;

// ----- Output vectors checking flags -------
	reg [0:0] c_flag;

// ----- Error counter: Deposit an error for config_done signal is not raised at the beginning -----
	integer nb_error= 1;
// ----- Number of clock cycles in configuration phase: 528 -----
// ----- Begin configuration done signal generation -----
initial
	begin
		__config_done__[0] = 1'b0;
	end

// ----- End configuration done signal generation -----

// ----- Begin raw programming clock signal generation -----
initial
	begin
		__prog_clock___reg__[0] = 1'b0;
	end
always
	begin
		#5	__prog_clock___reg__[0] = ~__prog_clock___reg__[0];
	end

// ----- End raw programming clock signal generation -----

// ----- Actual programming clock is triggered only when __config_done__ and __prog_reset__ are disabled -----
	assign __prog_clock__[0] = __prog_clock___reg__[0] & (~__config_done__[0]) & (~__prog_reset__[0]);

// ----- Begin raw operating clock signal generation -----
initial
	begin
		__op_clock___reg__[0] = 1'b0;
	end
always wait(~__greset__)
	begin
		#0.6491494179	__op_clock___reg__[0] = ~__op_clock___reg__[0];
	end

// ----- End raw operating clock signal generation -----
// ----- Actual operating clock is triggered only when __config_done__ is enabled -----
	assign __op_clock__[0] = __op_clock___reg__[0] & __config_done__[0];

// ----- Begin programming reset signal generation -----
initial
	begin
		__prog_reset__[0] = 1'b1;
	#10	__prog_reset__[0] = 1'b0;
	end

// ----- End programming reset signal generation -----

// ----- Begin programming set signal generation -----
initial
	begin
		__prog_set_[0] = 1'b1;
	#10	__prog_set_[0] = 1'b0;
	end

// ----- End programming set signal generation -----

// ----- Begin operating reset signal generation -----
// ----- Reset signal is enabled until the first clock cycle in operation phase -----
initial
	begin
		__greset__[0] = 1'b1;
	wait(__config_done__)
	#1.298298836	__greset__[0] = 1'b1;
	#2.596597672	__greset__[0] = 1'b0;
	end

// ----- End operating reset signal generation -----
// ----- Begin operating set signal generation: always disabled -----
initial
	begin
		__gset__[0] = 1'b0;
	end

// ----- End operating set signal generation: always disabled -----

// ----- Begin connecting global ports of FPGA fabric to stimuli -----
	assign clk[0] = __op_clock__[0];
	assign prog_clk[0] = __prog_clock__[0];
	assign reset[0] = __greset__[0];
	assign set[0] = __gset__[0];
// ----- End connecting global ports of FPGA fabric to stimuli -----
// ----- FPGA top-level module to be capsulated -----
	fpga_top FPGA_DUT (
		.prog_clk(prog_clk[0]),
		.set(set[0]),
		.reset(reset[0]),
		.clk(clk[0]),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[0:31]),
		.ccff_head(ccff_head[0]),
		.ccff_tail(ccff_tail[0]));

// ----- Link BLIF Benchmark I/Os to FPGA I/Os -----
// ----- Blif Benchmark input a is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD[6] -----
	assign gfpga_pad_GPIO_PAD[6] = a_shared_input[0];

// ----- Blif Benchmark input b is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD[17] -----
	assign gfpga_pad_GPIO_PAD[17] = b_shared_input[0];

// ----- Blif Benchmark output c is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD[4] -----
	assign c_fpga[0] = gfpga_pad_GPIO_PAD[4];

// ----- Wire unused FPGA I/Os to constants -----
	assign gfpga_pad_GPIO_PAD[0] = 1'b0;
	assign gfpga_pad_GPIO_PAD[1] = 1'b0;
	assign gfpga_pad_GPIO_PAD[2] = 1'b0;
	assign gfpga_pad_GPIO_PAD[3] = 1'b0;
	assign gfpga_pad_GPIO_PAD[5] = 1'b0;
	assign gfpga_pad_GPIO_PAD[7] = 1'b0;
	assign gfpga_pad_GPIO_PAD[8] = 1'b0;
	assign gfpga_pad_GPIO_PAD[9] = 1'b0;
	assign gfpga_pad_GPIO_PAD[10] = 1'b0;
	assign gfpga_pad_GPIO_PAD[11] = 1'b0;
	assign gfpga_pad_GPIO_PAD[12] = 1'b0;
	assign gfpga_pad_GPIO_PAD[13] = 1'b0;
	assign gfpga_pad_GPIO_PAD[14] = 1'b0;
	assign gfpga_pad_GPIO_PAD[15] = 1'b0;
	assign gfpga_pad_GPIO_PAD[16] = 1'b0;
	assign gfpga_pad_GPIO_PAD[18] = 1'b0;
	assign gfpga_pad_GPIO_PAD[19] = 1'b0;
	assign gfpga_pad_GPIO_PAD[20] = 1'b0;
	assign gfpga_pad_GPIO_PAD[21] = 1'b0;
	assign gfpga_pad_GPIO_PAD[22] = 1'b0;
	assign gfpga_pad_GPIO_PAD[23] = 1'b0;
	assign gfpga_pad_GPIO_PAD[24] = 1'b0;
	assign gfpga_pad_GPIO_PAD[25] = 1'b0;
	assign gfpga_pad_GPIO_PAD[26] = 1'b0;
	assign gfpga_pad_GPIO_PAD[27] = 1'b0;
	assign gfpga_pad_GPIO_PAD[28] = 1'b0;
	assign gfpga_pad_GPIO_PAD[29] = 1'b0;
	assign gfpga_pad_GPIO_PAD[30] = 1'b0;
	assign gfpga_pad_GPIO_PAD[31] = 1'b0;

// ----- Reference Benchmark Instanication -------
	or2 REF_DUT(
		.a(a_shared_input),
		.b(b_shared_input),
		.c(c_benchmark)
	);
// ----- End reference Benchmark Instanication -------

// ----- Begin bitstream loading during configuration phase -----
`define BITSTREAM_LENGTH 527
`define BITSTREAM_WIDTH 1
// ----- Virtual memory to store the bitstream from external file -----
reg [0:`BITSTREAM_WIDTH - 1] bit_mem[0:`BITSTREAM_LENGTH - 1];
reg [$clog2(`BITSTREAM_LENGTH):0] bit_index;
// ----- Registers used for fast configuration logic -----
reg [$clog2(`BITSTREAM_LENGTH):0] ibit;
reg [0:0] skip_bits;
// ----- Preload bitstream file to a virtual memory -----
initial begin
	$readmemb("fabric_bitstream.bit", bit_mem);
// ----- Configuration chain default input -----
	ccff_head[0] <= 1'b0;
	bit_index <= 0;
	skip_bits[0] <= 1'b0;
	for (ibit = 0; ibit < `BITSTREAM_LENGTH + 1; ibit = ibit + 1) begin
		if (1'b0 == bit_mem[ibit]) begin
			if (1'b1 == skip_bits[0]) begin
				bit_index <= bit_index + 1;
			end
		end else begin
			skip_bits[0] <= 1'b0;
		end
	end
end
// ----- 'else if' condition is required by Modelsim to synthesis the Verilog correctly -----
always @(negedge __prog_clock___reg__[0]) begin
	if (bit_index >= `BITSTREAM_LENGTH) begin
		__config_done__[0] <= 1'b1;
	end else if (bit_index >= 0 && bit_index < `BITSTREAM_LENGTH) begin
		ccff_head[0] <= bit_mem[bit_index];
		bit_index <= bit_index + 1;
	end
end
// ----- End bitstream loading during configuration phase -----

// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mux_ble4_out_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_4_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_4_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_5_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_5_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_6_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_6_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l3_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l3_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l4_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l4_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_4_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_4_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_5_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_5_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_6_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_6_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l3_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l3_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l4_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l4_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_4_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_4_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_5_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_5_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_6_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_6_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l3_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l3_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l4_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l4_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_4_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_4_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_5_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_5_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_6_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_6_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l3_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l3_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l4_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l4_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_4_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_4_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_5_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_5_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_6_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_6_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l3_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l3_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l4_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l4_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_4_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_4_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_5_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_5_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_6_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_6_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l3_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l3_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l4_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l4_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_4_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_4_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_5_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_5_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_6_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_6_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l3_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l3_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l4_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l4_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_4_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_4_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_5_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_5_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_6_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_6_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l3_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l3_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l4_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l4_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_4_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_4_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_5_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_5_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_6_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_6_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l3_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l3_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l4_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l4_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_4_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_4_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_5_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_5_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_6_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_6_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l3_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l3_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l4_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l4_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_4_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_4_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_5_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_5_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_6_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_6_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l3_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l3_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l4_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l4_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_4_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_4_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_5_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_5_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_6_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_6_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l3_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l3_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l4_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l4_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_4_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_4_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_5_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_5_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_6_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_6_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l3_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l3_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l4_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l4_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_4_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_4_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_5_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_5_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_6_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_6_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l3_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l3_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l4_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l4_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_4_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_4_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_5_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_5_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_6_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_6_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l3_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l3_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l4_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l4_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_4_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_4_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_5_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_5_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_6_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_6_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_3_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_3_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l3_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l3_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l4_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l4_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_0.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_0.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_0.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_0.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_12.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_12.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_12.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_12.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_12.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_12.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_12.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_12.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_0.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_0.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_0.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_0.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_2.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_2.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_2.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_2.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_2.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_2.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_2.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_2.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_12.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_12.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_12.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_12.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_12.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_12.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_12.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_12.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_14.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_14.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_14.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_14.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_14.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_14.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_14.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_14.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_2.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_2.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_2.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_2.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_2.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_2.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_4.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_4.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_4.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_4.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_4.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_4.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_6.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_6.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_6.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_6.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_6.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_6.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_8.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_8.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_8.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_8.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_8.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_8.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_10.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_10.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_10.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_10.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_10.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_10.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_14.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_14.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_14.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_14.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_14.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_14.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_16.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_16.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_16.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_16.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_16.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_16.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_24.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_24.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_24.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_24.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_24.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_24.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_4.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_4.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_4.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_4.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_4.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_4.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_6.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_6.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_6.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_6.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_6.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_6.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_8.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_8.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_8.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_8.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_8.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_8.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_10.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_10.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_10.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_10.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_10.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_10.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_16.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_16.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_16.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_16.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_16.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_16.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_24.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_24.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_24.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_24.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_24.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_24.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_18.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_18.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_18.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_18.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_20.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_20.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_20.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_20.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_22.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_22.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_22.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_top_track_22.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_18.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_18.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_18.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_18.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_20.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_20.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_20.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_20.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_22.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_22.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_22.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__0_.mux_right_track_22.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_0.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_0.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_0.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_0.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_12.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_12.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_12.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_12.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_12.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_12.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_12.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_12.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_1.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_1.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_1.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_1.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_3.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_3.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_3.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_3.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_15.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_15.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_15.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_15.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_2.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_2.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_2.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_2.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_2.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_2.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_4.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_4.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_4.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_4.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_4.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_4.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_6.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_6.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_6.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_6.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_6.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_6.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_8.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_8.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_8.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_8.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_8.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_8.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_10.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_10.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_10.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_10.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_10.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_10.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_14.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_14.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_14.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_14.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_14.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_14.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_16.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_16.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_16.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_16.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_16.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_16.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_24.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_24.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_24.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_24.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_24.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_24.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_5.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_5.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_7.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_7.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_11.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_11.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_13.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_13.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_18.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_18.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_18.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_18.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_20.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_20.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_20.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_20.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_22.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_22.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_22.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_right_track_22.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_19.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_19.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_19.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_19.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_21.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_21.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_21.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_21.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_23.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_23.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_23.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_23.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_25.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_25.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_25.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_0__1_.mux_bottom_track_25.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_0.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_0.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_0.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_0.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_2.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_2.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_2.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_2.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_2.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_2.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_2.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_2.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_14.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_14.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_14.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_14.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_14.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_14.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_14.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_14.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_1.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_1.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_1.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_1.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_3.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_3.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_3.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_3.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_3.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_3.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_3.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_3.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_13.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_13.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_13.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_13.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_13.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_13.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_13.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_13.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_15.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_15.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_15.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_15.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_15.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_15.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_15.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_15.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_4.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_4.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_4.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_4.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_4.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_4.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_6.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_6.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_6.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_6.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_6.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_6.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_8.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_8.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_8.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_8.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_8.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_8.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_10.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_10.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_10.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_10.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_10.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_10.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_12.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_12.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_12.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_12.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_12.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_12.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_16.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_16.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_16.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_16.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_16.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_16.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_5.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_5.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_5.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_5.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_5.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_5.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_7.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_7.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_7.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_7.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_7.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_7.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_9.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_9.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_9.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_9.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_9.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_9.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_11.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_11.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_11.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_11.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_11.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_11.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_17.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_17.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_17.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_17.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_17.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_17.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_25.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_25.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_25.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_25.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_25.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_25.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_18.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_18.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_18.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_18.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_20.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_20.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_20.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_20.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_22.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_22.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_22.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_22.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_24.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_24.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_24.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_top_track_24.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_19.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_19.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_19.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_19.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_21.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_21.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_21.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_21.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_23.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_23.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_23.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__0_.mux_left_track_23.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_1.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_1.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_1.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_1.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_13.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_13.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_13.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_13.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_1.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_1.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_1.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_1.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_13.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_13.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_13.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_13.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_13.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_13.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_13.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_13.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_3.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_3.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_5.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_5.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_7.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_7.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_11.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_11.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_15.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_15.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_25.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_25.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_25.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_25.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_25.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_25.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_3.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_3.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_3.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_3.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_3.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_3.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_5.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_5.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_5.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_5.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_5.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_5.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_7.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_7.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_7.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_7.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_7.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_7.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_9.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_9.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_9.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_9.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_9.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_9.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_11.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_11.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_11.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_11.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_11.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_11.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_15.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_15.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_15.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_15.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_15.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_15.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_17.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_17.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_17.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_17.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_17.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_17.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_25.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_25.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_25.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_25.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_25.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_25.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_19.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_19.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_19.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_19.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_21.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_21.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_21.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_21.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_23.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_23.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_23.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_bottom_track_23.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_19.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_19.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_19.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_19.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_21.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_21.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_21.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_21.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_23.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_23.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_23.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.sb_1__1_.mux_left_track_23.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_0.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_1.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_1.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_2.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_2.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_2.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_2.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_2.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_bottom_ipin_2.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_0.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_0.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_0.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_0.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_0.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_0.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_1.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_1.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_1.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_1.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_1.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_1.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_2.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_2.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_2.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_2.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_2.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_2.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_3.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_3.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_3.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_3.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_3.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_3.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_3.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_3.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_3.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_4.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_4.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_4.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_4.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_4.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_4.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_4.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_4.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_4.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_5.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_5.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_5.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_5.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_5.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_5.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_5.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_5.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_5.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_6.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_6.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_6.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_6.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_6.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_6.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_6.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_6.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_6.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_6.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_7.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_7.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_7.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_7.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_7.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_7.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__0_.mux_top_ipin_7.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_0.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_0.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_0.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_0.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_1.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_1.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_2.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_2.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_2.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_2.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_3.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_3.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_3.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_3.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_4.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_4.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_4.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_4.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_5.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_5.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_5.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_5.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_6.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_6.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_6.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_6.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_7.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_7.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_7.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_bottom_ipin_7.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_0.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_0.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_0.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_0.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_0.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_1.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_1.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_1.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_1.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_1.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_1.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_2.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_2.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_2.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_2.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_2.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cbx_1__1_.mux_top_ipin_2.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_0.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_0.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_0.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_0.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_0.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_1.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_1.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_1.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_1.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_1.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_1.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_left_ipin_1.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_0.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_0.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_0.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_0.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_0.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_0.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_1.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_1.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_1.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_1.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_1.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_1.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_2.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_2.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_2.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_2.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_2.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_2.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_3.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_3.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_3.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_3.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_3.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_3.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_3.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_3.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_4.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_4.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_4.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_4.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_4.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_4.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_4.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_4.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_4.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_5.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_5.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_5.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_5.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_5.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_5.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_5.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_6.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_6.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_6.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_6.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_6.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_6.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_6.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_6.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_6.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_7.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_7.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_7.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_7.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_7.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_7.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_7.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_7.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_0__1_.mux_right_ipin_7.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_0.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_0.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_0.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_0.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_0.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_1.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_1.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_1.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_1.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_1.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_1.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_1.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_2.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_2.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_2.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_2.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_2.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_2.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_2.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_2.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_2.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_2.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_2.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_2.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_3.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_3.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_3.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_3.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_3.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_3.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_3.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_3.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_3.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_3.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_3.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_4.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_4.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_4.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_4.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_4.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_4.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_4.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_4.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_4.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_4.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_4.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_4.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_5.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_5.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_5.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_5.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_5.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_5.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_5.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_5.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_5.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_5.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_5.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_5.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_6.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_6.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_6.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_6.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_6.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_6.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_6.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_6.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_6.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_6.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_6.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_6.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_7.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_7.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_7.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_7.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_7.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_7.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_7.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_7.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_7.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_7.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_7.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_left_ipin_7.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_0.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_0.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_0.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_0.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_0.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_0.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_1.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_1.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_1.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_1.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_1.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_1.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_2.mux_l1_in_2_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_2.mux_l1_in_2_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_2.mux_l2_in_1_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_2.mux_l2_in_1_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_2.mux_l3_in_0_.TGATE_0_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ------ BEGIN driver initialization -----
	initial begin
		$deposit(FPGA_DUT.cby_1__1_.mux_right_ipin_2.mux_l3_in_0_.TGATE_1_.in, $random % 2 ? 1'b1 : 1'b0);
	end
// ------ END driver initialization -----
// ----- Begin reset signal generation -----
// ----- Input Initialization -------
	initial begin
		a_shared_input <= 1'b0;
		b_shared_input <= 1'b0;

		c_flag[0] <= 1'b0;
	end

// ----- Input Stimulus -------
	always@(negedge __op_clock__[0]) begin
		a_shared_input <= $random;
		b_shared_input <= $random;
	end

// ----- Begin checking output vectors -------
// ----- Skip the first falling edge of clock, it is for initialization -------
	reg [0:0] sim_start;

	always@(negedge __op_clock__[0]) begin
		if (1'b1 == sim_start[0]) begin
			sim_start[0] <= ~sim_start[0];
		end else 
if (1'b1 == __config_done__) begin
			if(!(c_fpga === c_benchmark) && !(c_benchmark === 1'bx)) begin
				c_flag <= 1'b1;
			end else begin
				c_flag<= 1'b0;
			end
		end
	end

	always@(posedge c_flag) begin
		if(c_flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on c_fpga at time = %t", $realtime);
		end
	end


// ----- Configuration done must be raised in the end -------
	always@(posedge __config_done__[0]) begin
		nb_error = nb_error - 1;
	end

// ----- Begin output waveform to VCD file-------
	initial begin
		$dumpfile("or2_formal.vcd");
		$dumpvars(1, or2_autocheck_top_tb);
	end
// ----- END output waveform to VCD file -------

initial begin
	sim_start[0] <= 1'b1;
	$timeformat(-9, 2, "ns", 20);
	$display("Simulation start");
// ----- Can be changed by the user for his/her need -------
	#5312
	if(nb_error == 0) begin
		$display("Simulation Succeed");
	end else begin
		$display("Simulation Failed with %d error(s)", nb_error);
	end
	$finish;
end

endmodule
// ----- END Verilog module for or2_autocheck_top_tb -----

//----- Default net type -----
`default_nettype none

